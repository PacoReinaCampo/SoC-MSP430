// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/verunilibs/data/glbl.v,v 1.11 2005/03/15 02:06:36 nandinip Exp $

`timescale  1 ps / 1 ps

module glbl ();

  parameter ROC_WIDTH = 100000;
  parameter TOC_WIDTH = 0;

  wire GSR;
  wire GTS;
  wire PRLD;

  reg GSR_int;
  reg GTS_int;
  reg PRLD_int;

  //--------   JTAG Globals --------------
  wire JTAG_TDO_GLBL;
  wire JTAG_TCK_GLBL;
  wire JTAG_TDI_GLBL;
  wire JTAG_TMS_GLBL;
  wire JTAG_TRST_GLBL;

  reg JTAG_CAPTURE_GLBL;
  reg JTAG_RESET_GLBL;
  reg JTAG_SHIFT_GLBL;
  reg JTAG_UPDATE_GLBL;

  reg JTAG_SEL1_GLBL = 0;
  reg JTAG_SEL2_GLBL = 0 ;
  reg JTAG_SEL3_GLBL = 0;
  reg JTAG_SEL4_GLBL = 0;

  reg JTAG_USER_TDO1_GLBL = 1'bz;
  reg JTAG_USER_TDO2_GLBL = 1'bz;
  reg JTAG_USER_TDO3_GLBL = 1'bz;
  reg JTAG_USER_TDO4_GLBL = 1'bz;

  assign (weak1, weak0) GSR = GSR_int;
  assign (weak1, weak0) GTS = GTS_int;
  assign (weak1, weak0) PRLD = PRLD_int;

  initial begin
    GSR_int = 1'b1;
    PRLD_int = 1'b1;
    #(ROC_WIDTH)
    GSR_int = 1'b0;
    PRLD_int = 1'b0;
  end

  initial begin
    GTS_int = 1'b1;
    #(TOC_WIDTH)
    GTS_int = 1'b0;
  end

endmodule
