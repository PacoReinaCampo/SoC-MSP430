../../../../../bench/verilog/regression/leds.sv