////////////////////////////////////////////////////////////////////////////////
//                                            __ _      _     _               //
//                                           / _(_)    | |   | |              //
//                __ _ _   _  ___  ___ _ __ | |_ _  ___| | __| |              //
//               / _` | | | |/ _ \/ _ \ '_ \|  _| |/ _ \ |/ _` |              //
//              | (_| | |_| |  __/  __/ | | | | | |  __/ | (_| |              //
//               \__, |\__,_|\___|\___|_| |_|_| |_|\___|_|\__,_|              //
//                  | |                                                       //
//                  |_|                                                       //
//                                                                            //
//                                                                            //
//              MPSoC-MSP430 CPU                                              //
//              Multi Processor System on Chip                                //
//              BackBone Bus Interface                                       //
//                                                                            //
////////////////////////////////////////////////////////////////////////////////
// Copyright (c) 2019-2020 by the author(s)
//
// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
//
// The above copyright notice and this permission notice shall be included in
// all copies or substantial portions of the Software.
//
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
// THE SOFTWARE.
//
////////////////////////////////////////////////////////////////////////////////
// Author(s):
//   Paco Reina Campo <pacoreinacampo@queenfield.tech>

0 : bb_dout_o =  32'h1820e020;
1 : bb_dout_o =  32'ha8211000;
2 : bb_dout_o =  32'h1840e000;
3 : bb_dout_o =  32'h8462001c;
4 : bb_dout_o =  32'he4030000;
5 : bb_dout_o =  32'h10000000;
6 : bb_dout_o =  32'h15000000;
7 : bb_dout_o =  32'h84820020;
8 : bb_dout_o =  32'h9c400000;
9 : bb_dout_o =  32'hd4011000;
10 : bb_dout_o =  32'h9c600800;
11 : bb_dout_o =  32'hd4011804;
12 : bb_dout_o =  32'hd4012008;
13 : bb_dout_o =  32'hd401100c;
14 : bb_dout_o =  32'h9ca00001;
15 : bb_dout_o =  32'hd4012810;
16 : bb_dout_o =  32'hd4012814;
17 : bb_dout_o =  32'h84e10014;
18 : bb_dout_o =  32'hbc070001;
19 : bb_dout_o =  32'h0ffffffe;
20 : bb_dout_o =  32'h15000000;
21 : bb_dout_o =  32'h9c402000;
22 : bb_dout_o =  32'hd4011000;
23 : bb_dout_o =  32'h9c600800;
24 : bb_dout_o =  32'hd4011804;
25 : bb_dout_o =  32'h9c800001;
26 : bb_dout_o =  32'hd4012008;
27 : bb_dout_o =  32'hd401100c;
28 : bb_dout_o =  32'h9ca00001;
29 : bb_dout_o =  32'hd4012810;
30 : bb_dout_o =  32'hd4012814;
31 : bb_dout_o =  32'h84e10014;
32 : bb_dout_o =  32'hbc070001;
33 : bb_dout_o =  32'h0ffffffe;
34 : bb_dout_o =  32'h15000000;
35 : bb_dout_o =  32'h9c200100;
36 : bb_dout_o =  32'h44000800;
37 : bb_dout_o =  32'h15000000;
